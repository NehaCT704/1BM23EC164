package alu_pkg;

  typedef enum logic [1:0] {
    ADD,
    SUB,
    MUL,
    XOR
  } opcode_t;

endpackage
