// ----------------------------------------------------------------------------------
// File        : tb_traffic.sv
// Author      : Neha C T / 1BM23EC164
// Created     : 2026-02-04
// Module      : tb_traffic
// Project     : SystemVerilog and Verification (23EC6PE2SV),
//               Faculty: Prof. Ajaykumar Devarapalli
//
// Description : Simple testbench for Traffic Light Controller. Randomizes inputs and uses a 
//               covergroup to measure input combination coverage..
// ----------------------------------------------------------------------------------
